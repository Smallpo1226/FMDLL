
module FDE(Q,in,out);
input Q,w2;
output w1;
supply1 VDD;
supply0 VSS;
wire wire1,wire2;




endmodule