##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Mon Apr  1 12:10:47 2024
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO FMDLL
  CLASS BLOCK ;
  SIZE 72.800000 BY 70.560000 ;
  FOREIGN FMDLL 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN M[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8746 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.01339 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09 LAYER M2  ;
    ANTENNAMAXAREACAR 21.9022 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 0.156 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA2  ;
    ANTENNAMAXCUTCAR 0.375556 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 1.9068 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0139 LAYER M3  ;
    ANTENNAGATEAREA 0.241 LAYER M3  ;
    ANTENNAMAXAREACAR 40.4914 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 0.294502 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA3  ;
    ANTENNAMAXCUTCAR 0.874886 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.6594 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.00485 LAYER M4  ;
    ANTENNAGATEAREA 0.241 LAYER M4  ;
    ANTENNAMAXAREACAR 43.2275 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 0.314626 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA4  ;
    ANTENNAMAXCUTCAR 0.945011 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 1.953 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.01409 LAYER M5  ;
    ANTENNAGATEAREA 0.426 LAYER M5  ;
    ANTENNAMAXAREACAR 47.812 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 0.347701 LAYER M5  ;
    ANTENNAMAXCUTCAR 0.945011 LAYER VIA5  ;
    PORT
      LAYER M2 ;
        RECT 14.490000 70.060000 14.630000 70.560000 ;
    END
  END M[1]
  PIN M[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9275 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.006625 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.7378 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.00541 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.07 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.00064 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 8.1858 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.05861 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 2.8546 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 0.02053 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.059 LAYER M6  ;
    ANTENNAMAXAREACAR 55.4102 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 0.40839 LAYER M6  ;
    ANTENNAMAXCUTCAR 1.4322 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT -0.070000 70.060000 0.070000 70.560000 ;
    END
  END M[0]
  PIN N[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5747 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.004105 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 4.9714 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.03565 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 1.0906 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.00793 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.268 LAYER M4  ;
    ANTENNAMAXAREACAR 19.7241 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 0.143565 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.626393 LAYER VIA4  ;
    PORT
      LAYER M2 ;
        RECT 72.730000 70.060000 72.870000 70.560000 ;
    END
  END N[3]
  PIN N[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8319 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.013785 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.374 LAYER M2  ;
    ANTENNAMAXAREACAR 6.1703 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 0.0443583 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA2  ;
    ANTENNAMAXCUTCAR 0.237233 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.07 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.00064 LAYER M3  ;
    ANTENNAGATEAREA 0.374 LAYER M3  ;
    ANTENNAMAXAREACAR 6.35746 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 0.0460695 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA3  ;
    ANTENNAMAXCUTCAR 0.28242 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 2.2274 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.01605 LAYER M4  ;
    ANTENNAGATEAREA 0.374 LAYER M4  ;
    ANTENNAMAXAREACAR 12.3131 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 0.088984 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA4  ;
    ANTENNAMAXCUTCAR 0.327607 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.0714 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.00065 LAYER M5  ;
    ANTENNAGATEAREA 0.374 LAYER M5  ;
    ANTENNAMAXAREACAR 12.504 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 0.0907219 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA5  ;
    ANTENNAMAXCUTCAR 0.372794 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 2.5802 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 0.01857 LAYER M6  ;
    ANTENNAGATEAREA 0.514 LAYER M6  ;
    ANTENNAMAXAREACAR 17.5238 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 0.12685 LAYER M6  ;
    ANTENNAMAXCUTCAR 0.603571 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 58.170000 70.060000 58.310000 70.560000 ;
    END
  END N[2]
  PIN N[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8987 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.021265 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.282 LAYER M2  ;
    ANTENNAMAXAREACAR 11.5512 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 0.0829078 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA2  ;
    ANTENNAMAXCUTCAR 0.251975 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.07 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.00064 LAYER M3  ;
    ANTENNAGATEAREA 0.282 LAYER M3  ;
    ANTENNAMAXAREACAR 11.7995 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 0.0851773 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA3  ;
    ANTENNAMAXCUTCAR 0.311904 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 0.2282 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.00177 LAYER M4  ;
    ANTENNAGATEAREA 0.282 LAYER M4  ;
    ANTENNAMAXAREACAR 12.6087 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 0.0914539 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA4  ;
    ANTENNAMAXCUTCAR 0.371833 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.07 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.00064 LAYER M5  ;
    ANTENNAGATEAREA 0.282 LAYER M5  ;
    ANTENNAMAXAREACAR 12.8569 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 0.0937234 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA5  ;
    ANTENNAMAXCUTCAR 0.431762 LAYER VIA5  ;
    ANTENNAPARTIALMETALAREA 4.9322 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 0.03537 LAYER M6  ;
    ANTENNAGATEAREA 0.422 LAYER M6  ;
    ANTENNAMAXAREACAR 24.5446 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 0.177539 LAYER M6  ;
    ANTENNAMAXCUTCAR 0.603571 LAYER VIA6  ;
    PORT
      LAYER M2 ;
        RECT 43.610000 70.060000 43.750000 70.560000 ;
    END
  END N[1]
  PIN N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9508 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0285 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.563 LAYER M2  ;
    ANTENNAMAXAREACAR 8.96202 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 0.0652371 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA2  ;
    ANTENNAMAXCUTCAR 0.290018 LAYER VIA2  ;
    ANTENNAPARTIALMETALAREA 0.5418 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.00401 LAYER M3  ;
    ANTENNAGATEAREA 0.793 LAYER M3  ;
    ANTENNAMAXAREACAR 9.64525 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 0.0702938 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.375556 LAYER VIA3  ;
    PORT
      LAYER M2 ;
        RECT 29.050000 70.060000 29.190000 70.560000 ;
    END
  END N[0]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4371 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.010265 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.14 LAYER M3  ;
    ANTENNAMAXAREACAR 13.3346 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 0.0950714 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.241429 LAYER VIA3  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 35.210000 0.500000 35.350000 ;
    END
  END rst_n
  PIN clk_ext
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9275 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.006625 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 6.8922 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.04937 LAYER M4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.282 LAYER M4  ;
    ANTENNAMAXAREACAR 28.2521 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 0.208238 LAYER M4  ;
    ANTENNAMAXCUTCAR 0.845 LAYER VIA4  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 -0.070000 0.500000 0.070000 ;
    END
  END clk_ext
  PIN clk_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4947 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.032105 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 1.2082 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.00877 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA4  ;
    ANTENNAPARTIALMETALAREA 0.189 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.00149 LAYER M5  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA5  ;
    ANTENNADIFFAREA 0.322 LAYER M6  ;
    ANTENNAPARTIALMETALAREA 3.3642 LAYER M6  ;
    ANTENNAPARTIALMETALSIDEAREA 0.02417 LAYER M6  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.081 LAYER M6  ;
    ANTENNAMAXAREACAR 6.77663 LAYER M6  ;
    ANTENNAMAXSIDEAREACAR 0.0495433 LAYER M6  ;
    ANTENNAMAXCUTCAR 0.141845 LAYER VIA6  ;
    PORT
      LAYER M3 ;
        RECT 72.300000 -0.070000 72.800000 0.070000 ;
    END
  END clk_out
  PIN Sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END Sel[1]
  PIN Sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3517 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.009795 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.546 LAYER M3  ;
    ANTENNAMAXAREACAR 5.19249 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 0.0380678 LAYER M3  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA3  ;
    ANTENNAMAXCUTCAR 0.12381 LAYER VIA3  ;
    ANTENNAPARTIALMETALAREA 3.4034 LAYER M4  ;
    ANTENNAPARTIALMETALSIDEAREA 0.02445 LAYER M4  ;
    ANTENNAGATEAREA 0.546 LAYER M4  ;
    ANTENNAMAXAREACAR 11.4258 LAYER M4  ;
    ANTENNAMAXSIDEAREACAR 0.082848 LAYER M4  ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA4  ;
    ANTENNAMAXCUTCAR 0.154762 LAYER VIA4  ;
    ANTENNADIFFAREA 0.322 LAYER M5  ;
    ANTENNAPARTIALMETALAREA 2.5802 LAYER M5  ;
    ANTENNAPARTIALMETALSIDEAREA 0.01857 LAYER M5  ;
    ANTENNAGATEAREA 0.546 LAYER M5  ;
    ANTENNAMAXAREACAR 16.1515 LAYER M5  ;
    ANTENNAMAXSIDEAREACAR 0.116859 LAYER M5  ;
    ANTENNAMAXCUTCAR 0.154762 LAYER VIA5  ;
    PORT
      LAYER M3 ;
        RECT 0.000000 70.490000 0.500000 70.630000 ;
    END
  END Sel[0]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 70.800000 65.790000 72.800000 67.790000 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000000 65.790000 2.000000 67.790000 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.800000 2.770000 72.800000 4.770000 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000000 2.770000 2.000000 4.770000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.030000 68.560000 70.030000 70.560000 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.030000 0.000000 70.030000 2.000000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.770000 68.560000 4.770000 70.560000 ;
    END
    PORT
      LAYER M4 ;
        RECT 2.770000 0.000000 4.770000 2.000000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 70.800000 68.290000 72.800000 70.290000 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000000 68.290000 2.000000 70.290000 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.800000 0.270000 72.800000 2.270000 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000000 0.270000 2.000000 2.270000 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.530000 68.560000 72.530000 70.560000 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.530000 0.000000 72.530000 2.000000 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.270000 68.560000 2.270000 70.560000 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.270000 0.000000 2.270000 2.000000 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 72.800000 70.560000 ;
    LAYER M2 ;
      RECT 59.810000 68.560000 71.230000 70.560000 ;
      RECT 45.250000 68.560000 56.670000 70.560000 ;
      RECT 30.690000 68.560000 42.110000 70.560000 ;
      RECT 16.130000 68.560000 27.550000 70.560000 ;
      RECT 1.570000 68.560000 12.990000 70.560000 ;
      RECT 0.000000 0.000000 72.800000 68.560000 ;
    LAYER M3 ;
      RECT 2.000000 68.990000 72.800000 70.560000 ;
      RECT 0.000000 36.850000 72.800000 68.990000 ;
      RECT 2.000000 33.710000 72.800000 36.850000 ;
      RECT 0.000000 1.570000 72.800000 33.710000 ;
      RECT 2.000000 0.000000 70.800000 1.570000 ;
    LAYER M4 ;
      RECT 6.270000 67.060000 66.530000 70.560000 ;
      RECT 0.000000 3.500000 72.800000 67.060000 ;
      RECT 6.270000 0.000000 66.530000 3.500000 ;
    LAYER M5 ;
      RECT 3.500000 64.290000 69.300000 70.560000 ;
      RECT 0.000000 6.270000 72.800000 64.290000 ;
      RECT 3.500000 0.000000 69.300000 6.270000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 72.800000 70.560000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 72.800000 70.560000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 72.800000 70.560000 ;
  END
END FMDLL

END LIBRARY
