module FD_M( rst_n , M , DIV_m , CLK_exit );
    reg [1:0]cnt_tmp;
    reg clk_tmp;
    reg [1:0]cnt;
	input [1:0]M;
	input rst_n;
    input CLK_exit;
	output reg DIV_m;


endmodule