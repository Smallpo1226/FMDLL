module FDL (
    input clk_in;
    input [5:0] Q;
    input [5:0] Qb;
    output clk_out;
);

endmodule