module FD_M( rst_n , N , DIV_N , CLK_out );
    reg [2:0]cnt_tmp;
    reg clk_tmp;
    reg [2:0]cnt;
	input [2:0]N;
	input rst_n;
    input CLK_out;
	output reg DIV_N;


endmodule